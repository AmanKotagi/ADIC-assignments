module and_gate(a,b,y);
input a,b;
output y;
and i1(y,a,b);
endmodule

